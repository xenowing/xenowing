//
// User core top-level
//
// Instantiated by the real top-level: apf_top
//

`default_nettype none

module core_top (

//
// physical connections
//

///////////////////////////////////////////////////
// clock inputs 74.25mhz. not phase aligned, so treat these domains as asynchronous

input   wire            clk_74a, // mainclk1
input   wire            clk_74b, // mainclk1 

///////////////////////////////////////////////////
// cartridge interface
// switches between 3.3v and 5v mechanically
// output enable for multibit translators controlled by pic32

// GBA AD[15:8]
inout   wire    [7:0]   cart_tran_bank2,
output  wire            cart_tran_bank2_dir,

// GBA AD[7:0]
inout   wire    [7:0]   cart_tran_bank3,
output  wire            cart_tran_bank3_dir,

// GBA A[23:16]
inout   wire    [7:0]   cart_tran_bank1,
output  wire            cart_tran_bank1_dir,

// GBA [7] PHI#
// GBA [6] WR#
// GBA [5] RD#
// GBA [4] CS1#/CS#
//     [3:0] unwired
inout   wire    [7:4]   cart_tran_bank0,
output  wire            cart_tran_bank0_dir,

// GBA CS2#/RES#
inout   wire            cart_tran_pin30,
output  wire            cart_tran_pin30_dir,
// when GBC cart is inserted, this signal when low or weak will pull GBC /RES low with a special circuit
// the goal is that when unconfigured, the FPGA weak pullups won't interfere.
// thus, if GBC cart is inserted, FPGA must drive this high in order to let the level translators
// and general IO drive this pin.
output  wire            cart_pin30_pwroff_reset,

// GBA IRQ/DRQ
inout   wire            cart_tran_pin31,
output  wire            cart_tran_pin31_dir,

// infrared
input   wire            port_ir_rx,
output  wire            port_ir_tx,
output  wire            port_ir_rx_disable, 

// GBA link port
inout   wire            port_tran_si,
output  wire            port_tran_si_dir,
inout   wire            port_tran_so,
output  wire            port_tran_so_dir,
inout   wire            port_tran_sck,
output  wire            port_tran_sck_dir,
inout   wire            port_tran_sd,
output  wire            port_tran_sd_dir,
 
///////////////////////////////////////////////////
// cellular psram 0 and 1, two chips (64mbit x2 dual die per chip)

output  wire    [21:16] cram0_a,
inout   wire    [15:0]  cram0_dq,
input   wire            cram0_wait,
output  wire            cram0_clk,
output  wire            cram0_adv_n,
output  wire            cram0_cre,
output  wire            cram0_ce0_n,
output  wire            cram0_ce1_n,
output  wire            cram0_oe_n,
output  wire            cram0_we_n,
output  wire            cram0_ub_n,
output  wire            cram0_lb_n,

output  wire    [21:16] cram1_a,
inout   wire    [15:0]  cram1_dq,
input   wire            cram1_wait,
output  wire            cram1_clk,
output  wire            cram1_adv_n,
output  wire            cram1_cre,
output  wire            cram1_ce0_n,
output  wire            cram1_ce1_n,
output  wire            cram1_oe_n,
output  wire            cram1_we_n,
output  wire            cram1_ub_n,
output  wire            cram1_lb_n,

///////////////////////////////////////////////////
// sdram, 512mbit 16bit

output  wire    [12:0]  dram_a,
output  wire    [1:0]   dram_ba,
inout   wire    [15:0]  dram_dq,
output  wire    [1:0]   dram_dqm,
output  wire            dram_clk,
output  wire            dram_cke,
output  wire            dram_ras_n,
output  wire            dram_cas_n,
output  wire            dram_we_n,

///////////////////////////////////////////////////
// sram, 1mbit 16bit

output  wire    [16:0]  sram_a,
inout   wire    [15:0]  sram_dq,
output  wire            sram_oe_n,
output  wire            sram_we_n,
output  wire            sram_ub_n,
output  wire            sram_lb_n,

///////////////////////////////////////////////////
// vblank driven by dock for sync in a certain mode

input   wire            vblank,

///////////////////////////////////////////////////
// i/o to 6515D breakout usb uart

output  wire            dbg_tx,
input   wire            dbg_rx,

///////////////////////////////////////////////////
// i/o pads near jtag connector user can solder to

output  wire            user1,
input   wire            user2,

///////////////////////////////////////////////////
// RFU internal i2c bus 

inout   wire            aux_sda,
output  wire            aux_scl,

///////////////////////////////////////////////////
// RFU, do not use
output  wire            vpll_feed,


//
// logical connections
//

///////////////////////////////////////////////////
// video, audio output to scaler
output  wire    [23:0]  video_rgb,
output  wire            video_rgb_clock,
output  wire            video_rgb_clock_90,
output  wire            video_de,
output  wire            video_skip,
output  wire            video_vs,
output  wire            video_hs,
    
output  wire            audio_mclk,
input   wire            audio_adc,
output  wire            audio_dac,
output  wire            audio_lrck,

///////////////////////////////////////////////////
// bridge bus connection
// synchronous to clk_74a
output  wire            bridge_endian_little,
input   wire    [31:0]  bridge_addr,
input   wire            bridge_rd,
output  reg     [31:0]  bridge_rd_data,
input   wire            bridge_wr,
input   wire    [31:0]  bridge_wr_data,

///////////////////////////////////////////////////
// controller data
// 
// key bitmap:
//   [0]    dpad_up
//   [1]    dpad_down
//   [2]    dpad_left
//   [3]    dpad_right
//   [4]    face_a
//   [5]    face_b
//   [6]    face_x
//   [7]    face_y
//   [8]    trig_l1
//   [9]    trig_r1
//   [10]   trig_l2
//   [11]   trig_r2
//   [12]   trig_l3
//   [13]   trig_r3
//   [14]   face_select
//   [15]   face_start
//   [31:28] type
// joy values - unsigned
//   [ 7: 0] lstick_x
//   [15: 8] lstick_y
//   [23:16] rstick_x
//   [31:24] rstick_y
// trigger values - unsigned
//   [ 7: 0] ltrig
//   [15: 8] rtrig
//
input   wire    [31:0]  cont1_key,
input   wire    [31:0]  cont2_key,
input   wire    [31:0]  cont3_key,
input   wire    [31:0]  cont4_key,
input   wire    [31:0]  cont1_joy,
input   wire    [31:0]  cont2_joy,
input   wire    [31:0]  cont3_joy,
input   wire    [31:0]  cont4_joy,
input   wire    [15:0]  cont1_trig,
input   wire    [15:0]  cont2_trig,
input   wire    [15:0]  cont3_trig,
input   wire    [15:0]  cont4_trig
    
);

// not using the IR port, so turn off both the LED, and
// disable the receive circuit to save power
assign port_ir_tx = 0;
assign port_ir_rx_disable = 1;

// bridge endianness
assign bridge_endian_little = 0;

// cart is unused, so set all level translators accordingly
// directions are 0:IN, 1:OUT
assign cart_tran_bank3 = 8'hzz;
assign cart_tran_bank3_dir = 1'b0;
assign cart_tran_bank2 = 8'hzz;
assign cart_tran_bank2_dir = 1'b0;
assign cart_tran_bank1 = 8'hzz;
assign cart_tran_bank1_dir = 1'b0;
assign cart_tran_bank0 = 4'hf;
assign cart_tran_bank0_dir = 1'b1;
assign cart_tran_pin30 = 1'b0;      // reset or cs2, we let the hw control it by itself
assign cart_tran_pin30_dir = 1'bz;
assign cart_pin30_pwroff_reset = 1'b0;  // hardware can control this
assign cart_tran_pin31 = 1'bz;      // input
assign cart_tran_pin31_dir = 1'b0;  // input

// link port is unused, set to input only to be safe
// each bit may be bidirectional in some applications
assign port_tran_so = 1'bz;
assign port_tran_so_dir = 1'b0;     // SO is output only
assign port_tran_si = 1'bz;
assign port_tran_si_dir = 1'b0;     // SI is input only
assign port_tran_sck = 1'bz;
assign port_tran_sck_dir = 1'b0;    // clock direction can change
assign port_tran_sd = 1'bz;
assign port_tran_sd_dir = 1'b0;     // SD is input and not used

// tie off the rest of the pins we are not using
assign cram0_a = 'h0;
assign cram0_dq = {16{1'bZ}};
assign cram0_clk = 0;
assign cram0_adv_n = 1;
assign cram0_cre = 0;
assign cram0_ce0_n = 1;
assign cram0_ce1_n = 1;
assign cram0_oe_n = 1;
assign cram0_we_n = 1;
assign cram0_ub_n = 1;
assign cram0_lb_n = 1;

assign cram1_a = 'h0;
assign cram1_dq = {16{1'bZ}};
assign cram1_clk = 0;
assign cram1_adv_n = 1;
assign cram1_cre = 0;
assign cram1_ce0_n = 1;
assign cram1_ce1_n = 1;
assign cram1_oe_n = 1;
assign cram1_we_n = 1;
assign cram1_ub_n = 1;
assign cram1_lb_n = 1;

assign dram_a = 'h0;
assign dram_ba = 'h0;
assign dram_dq = {16{1'bZ}};
assign dram_dqm = 'h0;
assign dram_clk = 'h0;
assign dram_cke = 'h0;
assign dram_ras_n = 'h1;
assign dram_cas_n = 'h1;
assign dram_we_n = 'h1;

assign sram_a = 'h0;
assign sram_dq = {16{1'bZ}};
assign sram_oe_n  = 1;
assign sram_we_n  = 1;
assign sram_ub_n  = 1;
assign sram_lb_n  = 1;

assign dbg_tx = 1'bZ;
assign user1 = 1'bZ;
assign aux_scl = 1'bZ;
assign vpll_feed = 1'bZ;


// for bridge write data, we just broadcast it to all bus devices
// for bridge read data, we have to mux it
// add your own devices here
always @(*) begin
    casex(bridge_addr)
    default: begin
        bridge_rd_data <= 0;
    end
    32'h10xxxxxx: begin
        // example
        // bridge_rd_data <= example_device_data;
        bridge_rd_data <= 0;
    end
    32'hF8xxxxxx: begin
        bridge_rd_data <= cmd_bridge_rd_data;
    end
    endcase
end


//
// host/target command handler
//
    wire            clk_74a_reset_n;                // driven by host commands, can be used as core-wide reset
    wire    [31:0]  cmd_bridge_rd_data;
    
// bridge host commands
// synchronous to clk_74a
    wire            status_boot_done = pll_core_locked_s; 
    wire            status_setup_done = pll_core_locked_s; // rising edge triggers a target command
    wire            status_running = clk_74a_reset_n; // we are running as soon as reset_n goes high

    wire            dataslot_requestread;
    wire    [15:0]  dataslot_requestread_id;
    wire            dataslot_requestread_ack = 1;
    wire            dataslot_requestread_ok = 1;

    wire            dataslot_requestwrite;
    wire    [15:0]  dataslot_requestwrite_id;
    wire    [31:0]  dataslot_requestwrite_size;
    wire            dataslot_requestwrite_ack = 1;
    wire            dataslot_requestwrite_ok = 1;

    wire            dataslot_update;
    wire    [15:0]  dataslot_update_id;
    wire    [31:0]  dataslot_update_size;
    
    wire            dataslot_allcomplete;

    wire     [31:0] rtc_epoch_seconds;
    wire     [31:0] rtc_date_bcd;
    wire     [31:0] rtc_time_bcd;
    wire            rtc_valid;

    wire            savestate_supported;
    wire    [31:0]  savestate_addr;
    wire    [31:0]  savestate_size;
    wire    [31:0]  savestate_maxloadsize;

    wire            savestate_start;
    wire            savestate_start_ack;
    wire            savestate_start_busy;
    wire            savestate_start_ok;
    wire            savestate_start_err;

    wire            savestate_load;
    wire            savestate_load_ack;
    wire            savestate_load_busy;
    wire            savestate_load_ok;
    wire            savestate_load_err;
    
    wire            osnotify_inmenu;

// bridge target commands
// synchronous to clk_74a

    reg             target_dataslot_read;       
    reg             target_dataslot_write;
    reg             target_dataslot_getfile;    // require additional param/resp structs to be mapped
    reg             target_dataslot_openfile;   // require additional param/resp structs to be mapped
    
    wire            target_dataslot_ack;        
    wire            target_dataslot_done;
    wire    [2:0]   target_dataslot_err;

    reg     [15:0]  target_dataslot_id;
    reg     [31:0]  target_dataslot_slotoffset;
    reg     [31:0]  target_dataslot_bridgeaddr;
    reg     [31:0]  target_dataslot_length;
    
    wire    [31:0]  target_buffer_param_struct; // to be mapped/implemented when using some Target commands
    wire    [31:0]  target_buffer_resp_struct;  // to be mapped/implemented when using some Target commands
    
// bridge data slot access
// synchronous to clk_74a

    wire    [9:0]   datatable_addr;
    wire            datatable_wren;
    wire    [31:0]  datatable_data;
    wire    [31:0]  datatable_q;

core_bridge_cmd icb (

    .clk                ( clk_74a ),
    .reset_n            ( clk_74a_reset_n ),

    .bridge_endian_little   ( bridge_endian_little ),
    .bridge_addr            ( bridge_addr ),
    .bridge_rd              ( bridge_rd ),
    .bridge_rd_data         ( cmd_bridge_rd_data ),
    .bridge_wr              ( bridge_wr ),
    .bridge_wr_data         ( bridge_wr_data ),
    
    .status_boot_done       ( status_boot_done ),
    .status_setup_done      ( status_setup_done ),
    .status_running         ( status_running ),

    .dataslot_requestread       ( dataslot_requestread ),
    .dataslot_requestread_id    ( dataslot_requestread_id ),
    .dataslot_requestread_ack   ( dataslot_requestread_ack ),
    .dataslot_requestread_ok    ( dataslot_requestread_ok ),

    .dataslot_requestwrite      ( dataslot_requestwrite ),
    .dataslot_requestwrite_id   ( dataslot_requestwrite_id ),
    .dataslot_requestwrite_size ( dataslot_requestwrite_size ),
    .dataslot_requestwrite_ack  ( dataslot_requestwrite_ack ),
    .dataslot_requestwrite_ok   ( dataslot_requestwrite_ok ),

    .dataslot_update            ( dataslot_update ),
    .dataslot_update_id         ( dataslot_update_id ),
    .dataslot_update_size       ( dataslot_update_size ),
    
    .dataslot_allcomplete   ( dataslot_allcomplete ),

    .rtc_epoch_seconds      ( rtc_epoch_seconds ),
    .rtc_date_bcd           ( rtc_date_bcd ),
    .rtc_time_bcd           ( rtc_time_bcd ),
    .rtc_valid              ( rtc_valid ),
    
    .savestate_supported    ( savestate_supported ),
    .savestate_addr         ( savestate_addr ),
    .savestate_size         ( savestate_size ),
    .savestate_maxloadsize  ( savestate_maxloadsize ),

    .savestate_start        ( savestate_start ),
    .savestate_start_ack    ( savestate_start_ack ),
    .savestate_start_busy   ( savestate_start_busy ),
    .savestate_start_ok     ( savestate_start_ok ),
    .savestate_start_err    ( savestate_start_err ),

    .savestate_load         ( savestate_load ),
    .savestate_load_ack     ( savestate_load_ack ),
    .savestate_load_busy    ( savestate_load_busy ),
    .savestate_load_ok      ( savestate_load_ok ),
    .savestate_load_err     ( savestate_load_err ),

    .osnotify_inmenu        ( osnotify_inmenu ),
    
    .target_dataslot_read       ( target_dataslot_read ),
    .target_dataslot_write      ( target_dataslot_write ),
    .target_dataslot_getfile    ( target_dataslot_getfile ),
    .target_dataslot_openfile   ( target_dataslot_openfile ),
    
    .target_dataslot_ack        ( target_dataslot_ack ),
    .target_dataslot_done       ( target_dataslot_done ),
    .target_dataslot_err        ( target_dataslot_err ),

    .target_dataslot_id         ( target_dataslot_id ),
    .target_dataslot_slotoffset ( target_dataslot_slotoffset ),
    .target_dataslot_bridgeaddr ( target_dataslot_bridgeaddr ),
    .target_dataslot_length     ( target_dataslot_length ),

    .target_buffer_param_struct ( target_buffer_param_struct ),
    .target_buffer_resp_struct  ( target_buffer_resp_struct ),
    
    .datatable_addr         ( datatable_addr ),
    .datatable_wren         ( datatable_wren ),
    .datatable_data         ( datatable_data ),
    .datatable_q            ( datatable_q )

);



////////////////////////////////////////////////////////////////////////////////////////



// video generation
// ~12,288,000 hz pixel clock
//
// we want our video mode of 320x240 @ 60hz, this results in 204800 clocks per frame
// we need to add hblank and vblank times to this, so there will be a nondisplay area. 
// it can be thought of as a border around the visible area.
// to make numbers simple, we can have 400 total clocks per line, and 320 visible.
// dividing 204800 by 400 results in 512 total lines per frame, and 240 visible.
// this pixel clock is fairly high for the relatively low resolution, but that's fine.
// PLL output has a minimum output frequency anyway.

// To ship video data from the system clock domain to the video output domain, we use a FIFO line buffer.
//  The line buffer is large enough to store two lines' worth of pixel data. While the line stored in the first
//   half is displayed, the following line's data can be written to the second half, and the halves are swapped
//   after each line.
//  When a vsync pulse is generated, both read and write pointers are reset to point to the beginning of the line
//   buffer.
//  When each line prior to a line which will be displayed begins, a pulse is generated and synchronized into the
//   system clock domain which triggers writing one line's worth of video data into the line buffer. The write
//   address is incremented modulo the full line buffer size after each pixel is written. Writes are disabled at
//   all other times.
//  For each pixel prior to a pixel which will be displayed on each line to be displayed, a read is issued to the
//   line buffer such that the pixel data will be ready on the following cycle when it will be displayed. The read
//   address is incremented modulo the full line buffer size after each pixel is read. Reads are disabled at all
//   other times.
//  As long as writing a line's worth of video data into the buffer always takes less time than reading/displaying
//   a line, the active read/write regions will never overlap, and all potential metastability errors are avoided.

    // Synchronize reset into video clock domain
    wire clk_core_12288_reset_n;
    SyncChain #(
        .STAGES(3)
    ) clk_core_12288_reset_n_sync_chain (
        .reset_n(clk_74a_reset_n),
        .clk(clk_core_12288),

        .x(clk_74a_reset_n),

        .x_sync(clk_core_12288_reset_n)
    );

assign video_rgb_clock = clk_core_12288;
assign video_rgb_clock_90 = clk_core_12288_90deg;
assign video_rgb = vidout_rgb;
assign video_de = vidout_de;
assign video_skip = vidout_skip;
assign video_vs = vidout_vs;
assign video_hs = vidout_hs;

    localparam  VID_V_BPORCH = 'd10;
    localparam  VID_V_ACTIVE = 'd240;
    localparam  VID_V_TOTAL = 'd512;
    localparam  VID_H_BPORCH = 'd10;
    localparam  VID_H_ACTIVE = 'd320;
    localparam  VID_H_TOTAL = 'd400;
    
    reg [9:0]   x_count;
    reg [9:0]   y_count;

    reg [23:0]  vidout_rgb;
    reg         vidout_de;
    reg         vidout_skip;
    reg         vidout_vs;
    reg         vidout_hs;

    reg vidout_write_line_pulse;

    reg video_line_buffer_read_enable;
    reg [9:0] video_line_buffer_read_addr;
    wire shovel_line_buffer_read_data;
    wire [23:0] test_pattern_line_buffer_read_data;

always @(posedge clk_core_12288 or negedge clk_core_12288_reset_n) begin

    if(~clk_core_12288_reset_n) begin
    
        x_count <= 0;
        y_count <= 0;

        vidout_write_line_pulse <= 1'b0;

        video_line_buffer_read_enable <= 1'b0;
        
    end else begin
        vidout_de <= 0;
        vidout_skip <= 0;
        vidout_vs <= 0;
        vidout_hs <= 0;
        
        // x and y counters
        x_count <= x_count + 1'b1;
        if(x_count == VID_H_TOTAL-1) begin
            x_count <= 0;
            
            y_count <= y_count + 1'b1;
            if(y_count == VID_V_TOTAL-1) begin
                y_count <= 0;
            end
        end
        
        // generate sync 
        if(x_count == 0 && y_count == 0) begin
            // sync signal in back porch
            // new frame
            vidout_vs <= 1;

            video_line_buffer_read_addr <= 10'd0;
        end
        
        // we want HS to occur a bit after VS, not on the same cycle
        if(x_count == 3) begin
            // sync signal in back porch
            // new line
            vidout_hs <= 1;
        end

        // issue line buffer write pulses
        //  These should occur on the beginning of every line that's prior to a line that will be displayed
        if (x_count == 0 && y_count >= VID_V_BPORCH - 1 && y_count < VID_V_ACTIVE+VID_V_BPORCH - 1) begin
            vidout_write_line_pulse <= 1'b1;
        end
        else begin
            vidout_write_line_pulse <= 1'b0;
        end

        // issue line buffer reads
        //  These need to occur one cycle before each displayed pixel
        video_line_buffer_read_enable <= 1'b0;
        if (y_count >= VID_V_BPORCH && y_count < VID_V_ACTIVE+VID_V_BPORCH) begin
            // Remember that we're setting up signals for the following cycle, so we offset x by 2 instead of 1.
            //  In other words, we want to issue reads a cycle early on the following cycle.
            if (x_count >= VID_H_BPORCH - 2 && x_count < VID_H_ACTIVE+VID_H_BPORCH - 2) begin
                video_line_buffer_read_enable <= 1'b1;
            end
        end
        // Next address should only increment if we actually performed a read this cycle
        if (video_line_buffer_read_enable) begin
            video_line_buffer_read_addr <= video_line_buffer_read_addr + 10'd1;
            if (video_line_buffer_read_addr == VID_H_ACTIVE * 2 - 1) begin
                video_line_buffer_read_addr <= 10'd0;
            end
        end

        // inactive screen areas are black
        vidout_rgb <= 24'h0;
        // generate active video
        if(x_count >= VID_H_BPORCH && x_count < VID_H_ACTIVE+VID_H_BPORCH) begin

            if(y_count >= VID_V_BPORCH && y_count < VID_V_ACTIVE+VID_V_BPORCH) begin
                // data enable. this is the active region of the line
                vidout_de <= 1;
                
                vidout_rgb <= shovel_line_buffer_read_data ? 24'hffffff : test_pattern_line_buffer_read_data;
                
            end 
        end
    end
end

    // Synchronize reset into sdram clock domain
    wire clk_sdram_reset_n;
    SyncChain #(
        .STAGES(3)
    ) clk_sdram_reset_n_sync_chain (
        .reset_n(clk_74a_reset_n),
        .clk(clk_sdram),

        .x(clk_74a_reset_n),

        .x_sync(clk_sdram_reset_n)
    );

    // Synchronize control pulses from video output domain to system domain
    wire system_write_vsync_pulse;
    CdcPulse p0 (
        .src_reset_n(clk_core_12288_reset_n),
        .src_clk(clk_core_12288),
        .src_pulse(vidout_vs),

        .dst_reset_n(clk_sdram_reset_n),
        .dst_clk(clk_sdram),
        .dst_pulse(system_write_vsync_pulse)
    );

    wire system_write_line_pulse;
    CdcPulse p1 (
        .src_reset_n(clk_core_12288_reset_n),
        .src_clk(clk_core_12288),
        .src_pulse(vidout_write_line_pulse),

        .dst_reset_n(clk_sdram_reset_n),
        .dst_clk(clk_sdram),
        .dst_pulse(system_write_line_pulse)
    );

    // Shovel line buffer
    wire shovel_line_buffer_write_enable;
    reg [9:0] shovel_line_buffer_write_addr;
    wire shovel_line_buffer_write_data;
    UnidirectionalDualPortBram #(
        .DATA(1),
        .ADDR(10),
        .DEPTH(VID_H_ACTIVE * 2)
    ) shovel_line_buffer (
        .write_clk(clk_sdram),
        .write_enable(shovel_line_buffer_write_enable),
        .write_addr(shovel_line_buffer_write_addr),
        .write_data(shovel_line_buffer_write_data),

        .read_clk(clk_core_12288),
        .read_enable(video_line_buffer_read_enable),
        .read_addr(video_line_buffer_read_addr),
        .read_data(shovel_line_buffer_read_data)
    );

    always @(posedge clk_sdram) begin
        if (system_write_vsync_pulse) begin
            shovel_line_buffer_write_addr <= 10'd0;
        end
        else if (shovel_line_buffer_write_enable) begin
            shovel_line_buffer_write_addr <= shovel_line_buffer_write_addr + 10'd1;
            if (shovel_line_buffer_write_addr == VID_H_ACTIVE * 2 - 1) begin
                shovel_line_buffer_write_addr <= 10'd0;
            end
        end
    end

    // Shovel
    // TODO: Figure out a good way to keep this consistent with kaze rtl
    localparam SHOVEL_BOOTLOADER_ADDR_BIT_WIDTH = 12;
    wire shovel_bootloader_bus_enable;
    wire [SHOVEL_BOOTLOADER_ADDR_BIT_WIDTH - 1:0] shovel_bootloader_bus_addr;
    wire shovel_bootloader_bus_write;
    wire [31:0] shovel_bootloader_bus_write_data;
    wire [3:0] shovel_bootloader_bus_write_byte_enable;
    wire [31:0] shovel_bootloader_bus_read_data;
    reg shovel_bootloader_bus_read_data_valid;
    Shovel shovel(
        .reset_n(clk_sdram_reset_n),
        .clk(clk_sdram),

        .system_write_vsync_pulse(system_write_vsync_pulse),
        .system_write_line_pulse(system_write_line_pulse),

        .video_line_buffer_write_enable(shovel_line_buffer_write_enable),
        .video_line_buffer_write_data(shovel_line_buffer_write_data),

        .bootloader_bus_ready(1'b1),
        .bootloader_bus_enable(shovel_bootloader_bus_enable),
        .bootloader_bus_addr(shovel_bootloader_bus_addr),
        .bootloader_bus_write(shovel_bootloader_bus_write),
        .bootloader_bus_write_data(shovel_bootloader_bus_write_data),
        .bootloader_bus_write_byte_enable(shovel_bootloader_bus_write_byte_enable),
        .bootloader_bus_read_data(shovel_bootloader_bus_read_data),
        .bootloader_bus_read_data_valid(shovel_bootloader_bus_read_data_valid)
    );

    always @(posedge clk_sdram) begin
        shovel_bootloader_bus_read_data_valid <= shovel_bootloader_bus_enable && !shovel_bootloader_bus_write;
    end

    // Test pattern line buffer
    wire test_pattern_line_buffer_write_enable;
    reg [9:0] test_pattern_line_buffer_write_addr;
    wire [23:0] test_pattern_line_buffer_write_data;
    UnidirectionalDualPortBram #(
        .DATA(24),
        .ADDR(10),
        .DEPTH(VID_H_ACTIVE * 2)
    ) test_pattern_line_buffer (
        .write_clk(clk_sdram),
        .write_enable(test_pattern_line_buffer_write_enable),
        .write_addr(test_pattern_line_buffer_write_addr),
        .write_data(test_pattern_line_buffer_write_data),

        .read_clk(clk_core_12288),
        .read_enable(video_line_buffer_read_enable),
        .read_addr(video_line_buffer_read_addr),
        .read_data(test_pattern_line_buffer_read_data)
    );

    always @(posedge clk_sdram) begin
        if (system_write_vsync_pulse) begin
            test_pattern_line_buffer_write_addr <= 10'd0;
        end
        else if (test_pattern_line_buffer_write_enable) begin
            test_pattern_line_buffer_write_addr <= test_pattern_line_buffer_write_addr + 10'd1;
            if (test_pattern_line_buffer_write_addr == VID_H_ACTIVE * 2 - 1) begin
                test_pattern_line_buffer_write_addr <= 10'd0;
            end
        end
    end

    // Test pattern generator
    VideoTestPatternGenerator test_pattern_generator(
        .reset_n(clk_sdram_reset_n),
        .clk(clk_sdram),

        .system_write_vsync_pulse(system_write_vsync_pulse),
        .system_write_line_pulse(system_write_line_pulse),

        .video_line_buffer_write_enable(test_pattern_line_buffer_write_enable),
        .video_line_buffer_write_data(test_pattern_line_buffer_write_data)
    );

    // Bootloader memory
    bootloader_mem shovel_bootloader_mem(
        .clock_a(clk_sdram),
        .address_a(shovel_bootloader_bus_addr),
        .rden_a(shovel_bootloader_bus_enable && !shovel_bootloader_bus_write),
        .wren_a(shovel_bootloader_bus_enable && shovel_bootloader_bus_write),
        .data_a(shovel_bootloader_bus_write_data),
        .byteena_a(shovel_bootloader_bus_write_byte_enable),
        .q_a(shovel_bootloader_bus_read_data),

        .clock_b(clk_74a),
        .address_b(bridge_addr[SHOVEL_BOOTLOADER_ADDR_BIT_WIDTH - 1 + 2:2]),
        .rden_b(1'b0),
        .wren_b(bridge_wr && bridge_addr[31:24] == 8'h10),
        // bridge_wr_data is big-endian
        .data_b({
            bridge_wr_data[7:0],
            bridge_wr_data[15:8],
            bridge_wr_data[23:16],
            bridge_wr_data[31:24]
        })
    );


//
// audio i2s silence generator
// see other examples for actual audio generation
//

assign audio_mclk = audgen_mclk;
assign audio_dac = audgen_dac;
assign audio_lrck = audgen_lrck;

// generate MCLK = 12.288mhz with fractional accumulator
    reg         [21:0]  audgen_accum;
    reg                 audgen_mclk;
    parameter   [20:0]  CYCLE_48KHZ = 21'd122880 * 2;
always @(posedge clk_74a) begin
    audgen_accum <= audgen_accum + CYCLE_48KHZ;
    if(audgen_accum >= 21'd742500) begin
        audgen_mclk <= ~audgen_mclk;
        audgen_accum <= audgen_accum - 21'd742500 + CYCLE_48KHZ;
    end
end

// generate SCLK = 3.072mhz by dividing MCLK by 4
    reg [1:0]   aud_mclk_divider;
    wire        audgen_sclk = aud_mclk_divider[1] /* synthesis keep*/;
    reg         audgen_lrck_1;
always @(posedge audgen_mclk) begin
    aud_mclk_divider <= aud_mclk_divider + 1'b1;
end

// shift out audio data as I2S 
// 32 total bits per channel, but only 16 active bits at the start and then 16 dummy bits
//
    reg     [4:0]   audgen_lrck_cnt;    
    reg             audgen_lrck;
    reg             audgen_dac;
always @(negedge audgen_sclk) begin
    audgen_dac <= 1'b0;
    // 48khz * 64
    audgen_lrck_cnt <= audgen_lrck_cnt + 1'b1;
    if(audgen_lrck_cnt == 31) begin
        // switch channels
        audgen_lrck <= ~audgen_lrck;
        
    end 
end


///////////////////////////////////////////////


    wire    clk_core_12288;
    wire    clk_core_12288_90deg;
    wire clk_sdram;
    
    wire    pll_core_locked;
    wire    pll_core_locked_s;
synch_3 s01(pll_core_locked, pll_core_locked_s, clk_74a);

mf_pllbase mp1 (
    .refclk         ( clk_74a ),
    .rst            ( 0 ),
    
    .outclk_0       ( clk_core_12288 ),
    .outclk_1       ( clk_core_12288_90deg ),
    .outclk_2(clk_sdram),
    
    .locked         ( pll_core_locked )
);


    
endmodule
