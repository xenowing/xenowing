`default_nettype none

module decode(
    input reset_n,
    input clk,

    output ready,
    input enable,

    input [31:0] instruction);

    // TODO

endmodule
