typedef enum [3:0] {
    ADD,
    SUB,
    AND,
    OR,
    XOR,
    SLL,
    SRL,
    SRA,
    EQ,
    NE,
    LT,
    LTU,
    GE,
    GEU
} alu_op_t;
